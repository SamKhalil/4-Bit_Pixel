*It should be included in the file you describe the circuit with:
*.lib photodiode.cir
*-----------------< Photo Diode Sub Ciruit >--------------------------------------------------
.SUBCKT PhotoDiode   N1_R1C1
.param  	Vsource = 5V
.param  	Ipd_1 = 200pA
VDD	 	VDD 	VSS 	DC     Vsource
VSS 		VSS 	0 	DC	 0
*----------The photodiode for Ith  PIXEL R1C1----------
I1_R1C1 	VDD	 	N1_R1C1 	 DC		Ipd_1
Mpd_R1C1	N1_R1C1 	N1_R1C1	 N1_R1C1	VDD	PM	W=10e-6 	L=0.6e-6
+ AD=50E-12 	PD=0 AS=50E-12 	PS=0

.ENDS	PhotoDiode   
*-----------------End Photo Diode---------------------------------------------------------
*Alternatively, add directly the following lines to your code
*I1_R1C1 VDD N1_R1C1 DC PHOTOCURRENT_R1C1
*Mpd_R1C1 N1_R1C1 N1_R1C1 N1_R1C1 VDD MP W=10e-6 L=0.6e-6 + AD=50E-12 PD=0 AS=50E-12 PS=0